module encoder (s0, s1, s2, s3, s4, s5, s6, in, enable);
	input enable;
	input [3:0] in;//declare as a 4bit binary
	output reg s0, s1, s2, s3, s4, s5, s6;

	always @(*) begin
	if(enable)begin
		if (in==4'b0000) begin
			s0=0;
			s1=0;
			s2=0;
			s3=0;
			s4=0;
			s5=0;
			s6=1;
		end
		else if (in==4'b0001) begin
			s0=1;
			s1=0;
			s2=0;
			s3=1;
			s4=1;
			s5=1;
			s6=1;
		end
		else if (in==4'b0010) begin
			s0=0;
			s1=0;
			s2=1;
			s3=0;
			s4=0;
			s5=1;
			s6=0;
		end
		else if (in==4'b0011) begin
			s0=0;
			s1=0;
			s2=0;
			s3=0;
			s4=1;
			s5=1;
			s6=0;
		end
		else if (in==4'b0100) begin
			s0=1;
			s1=0;
			s2=0;
			s3=1;
			s4=1;
			s5=0;
			s6=0;
		end
		else if (in==4'b0101) begin
			s0=0;
			s1=1;
			s2=0;
			s3=0;
			s4=1;
			s5=0;
			s6=0;
		end
		else if (in==4'b0110) begin
			s0=0;
			s1=1;
			s2=0;
			s3=0;
			s4=0;
			s5=0;
			s6=0;
		end
		else if (in==4'b0111) begin
			s0=0;
			s1=0;
			s2=0;
			s3=1;
			s4=1;
			s5=1;
			s6=1;
		end
		else if (in==4'b1000) begin
			s0=0;
			s1=0;
			s2=0;
			s3=0;
			s4=0;
			s5=0;
			s6=0;
		end
		else if (in==4'b1001) begin
			s0=0;
			s1=0;
			s2=0;
			s3=1;
			s4=1;
			s5=0;
			s6=0;
		end
		else if (in==4'b1010) begin
			s0=0;
			s1=0;
			s2=0;
			s3=1;
			s4=0;
			s5=0;
			s6=0;
		end
		else if (in==4'b1011) begin
			s0=1;
			s1=1;
			s2=0;
			s3=0;
			s4=0;
			s5=0;
			s6=0;
		end
		else if (in==4'b1100) begin
			s0=0;
			s1=1;
			s2=1;
			s3=0;
			s4=0;
			s5=0;
			s6=1;
		end
		else if (in==4'b1101) begin
			s0=1;
			s1=0;
			s2=0;
			s3=0;
			s4=0;
			s5=1;
			s6=0;
		end
		else if (in==4'b1110) begin
			s0=0;
			s1=1;
			s2=1;
			s3=0;
			s4=0;
			s5=0;
			s6=0;
		end
		else if (in==4'b1111) begin
			s0=0;
			s1=1;
			s2=1;
			s3=1;
			s4=0;
			s5=0;
			s6=0;
		end
		else begin
			s0=0;
			s1=0;
			s2=0;
			s3=1;
			s4=1;
			s5=1;
			s6=1;
		end
	end
	else begin
		s0 = 0;
		s1 = 0;
		s2 = 0;
		s3 = 0;
		s4 = 0;
		s5 = 0;
		s6 = 1;
	end
	end
endmodule 